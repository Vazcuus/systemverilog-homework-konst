//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module serial_to_parallel
# (
    parameter width = 8
)
(
    input                      clk,
    input                      rst,

    input                      serial_valid,
    input                      serial_data,

    output logic               parallel_valid,
    output logic [width - 1:0] parallel_data
);
    // Task:
    // Implement a module that converts single-bit serial data to the multi-bit parallel value.
    //
    // The module should accept one-bit values with valid interface in a serial manner.
    // After accumulating 'width' bits and receiving last 'serial_valid' input,
    // the module should assert the 'parallel_valid' at the same clock cycle
    // and output 'parallel_data' value.
    //
    // Note:
    // Check the waveform diagram in the README for better understanding.
    logic [2:0] bit_counter;

    logic [width - 1:0] data_reg;

    assign parallel_valid = (bit_counter == width - 1) && serial_valid;

    assign parallel_data = parallel_valid ? {serial_data, data_reg[width - 1:1]} : data_reg;

    always_ff @ (posedge clk, posedge rst)
        if (rst) begin
            bit_counter <= '0;
            data_reg    <= '0;
        end
        else 
        begin
        if (serial_valid) 
        begin
            data_reg <= {serial_data, data_reg[width - 1:1]};
            if (bit_counter == width - 1)
                bit_counter <= '0;
            else
                bit_counter <= bit_counter + 1;
        end
    end
endmodule
